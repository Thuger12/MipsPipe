module stageWB ();
endmodule 