module InstrMemory ();
endmodule 