module stageMem ();
endmodule 